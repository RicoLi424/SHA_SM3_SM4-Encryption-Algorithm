module SM3ProcessMessageBlock(clk,rst,enable,messageBlock,V_i,V_o);
    
	 //输入输出变量
    input  clk,rst,enable;          //输入变量：时钟，低电平有效异步复位信号，高电平有效使能信号
    input  [511:0] messageBlock;    //输入变量：压缩函数的输入变量之一B(i)，待处理消息块
	 input  [255:0] V_i;             //输入变量：压缩函数的输入变量之一V(i)，intermediate的旧值
    output [255:0] V_o;             //输出变量：压缩函数的输出变量V(i+1)，intermediate的新值
	 
    wire   clk,rst,enable;          //线网型
    wire   [511:0] messageBlock;    //线网型
	 wire   [255:0] V_i;             //线网型
	 reg    [255:0] V_o;             //寄存器型
	 
	 //中间变（常）量
    reg    [31:0]  Tj;              //常量Tj
	 reg    [5:0]   j;               //压缩次数
	 reg    [31:0]  A,B,C,D,E,F,G,H; //字寄存器，用于压缩
	 reg    [31:0]  SS1t;            //求中间变量SS1时所用的中间变量，为置换函数的自变量
	 reg    [31:0]  SS1,SS2,TT1,TT2; //压缩过程中的中间变量，暂存数据
	 reg    [31:0]  FF,GG;           //布尔函数
	 reg    [5:0]   count;           //消息扩展时所用的计数器
	 reg    [31:0]  w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15,
	                w16,w17,w18,w19,w20,w21,w22,w23,w24,w25,w26,w27,w28,w29,w30,w31,
	                w32,w33,w34,w35,w36,w37,w38,w39,w40,w41,w42,w43,w44,w45,w46,w47,
	                w48,w49,w50,w51,w52,w53,w54,w55,w56,w57,w58,w59,w60,w61,w62,w63,
	                w64,w65,w66,w67; //扩展后的部分消息，用于压缩时字寄存器内数据逻辑运算
						 
	 reg    [31:0]  w_0,w_1,w_2,w_3,w_4,w_5,w_6,w_7,w_8,w_9,w_10,w_11,w_12,w_13,w_14,w_15,
	                w_16,w_17,w_18,w_19,w_20,w_21,w_22,w_23,w_24,w_25,w_26,w_27,w_28,w_29,w_30,w_31,
	                w_32,w_33,w_34,w_35,w_36,w_37,w_38,w_39,w_40,w_41,w_42,w_43,w_44,w_45,w_46,w_47,
	                w_48,w_49,w_50,w_51,w_52,w_53,w_54,w_55,w_56,w_57,w_58,w_59,w_60,w_61,w_62,w_63;
						                  //扩展后的部分消息，用于压缩时字寄存器内数据逻辑运算
	 reg    [31:0]  wt_16,wt_17,wt_18,wt_19,wt_20,wt_21,wt_22,wt_23,wt_24,wt_25,wt_26,wt_27,wt_28,wt_29,wt_30,wt_31,
	                wt_32,wt_33,wt_34,wt_35,wt_36,wt_37,wt_38,wt_39,wt_40,wt_41,wt_42,wt_43,wt_44,wt_45,wt_46,wt_47,
	                wt_48,wt_49,wt_50,wt_51,wt_52,wt_53,wt_54,wt_55,wt_56,wt_57,wt_58,wt_59,wt_60,wt_61,wt_62,wt_63,
	                wt_64,wt_65,wt_66,wt_67;
	
	 
 
    //消息扩展部分
	 always@(posedge clk or negedge rst)
	 begin
	     if(!rst)
		  begin
		  //复位信号有效时，清零
		      count <= 6'd0;
		      {w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15} <= 256'd0;
		  end
		  else if(!enable)
		  begin
		  //使能信号无效时，停止工作
		      count <= count;
		  end
		  else
		  begin
		      case(count)
				    6'd0:
					 begin
					     {w0,w1,w2,w3,w4,w5,w6,w7,w8,w9,w10,w11,w12,w13,w14,w15} <= messageBlock;//计算w0-w15
						  
						  count <= count + 6'd1;//count自加一
					 end						  
					 6'd1:
					 begin    
					     wt_16 <= w0 ^ w7 ^ {w13[16:0],w13[31:17]};//中间变量
						  wt_17 <= w1 ^ w8 ^ {w14[16:0],w14[31:17]};
					     wt_18 <= w2 ^ w9 ^ {w15[16:0],w15[31:17]};
						  
						  w_0 <= w0 ^ w4;//计算w_0-w_11
						  w_1 <= w1 ^ w5;
						  w_2 <= w2 ^ w6;
						  w_3 <= w3 ^ w7;
						  w_4 <= w4 ^ w8;
						  w_5 <= w5 ^ w9;
						  w_6 <= w6 ^ w10;
						  w_7 <= w7 ^ w11;
						  w_8 <= w8 ^ w12;
						  w_9 <= w9 ^ w13;
						  w_10 <= w10 ^ w14;
						  w_11 <= w11 ^ w15;
						  
						  count <= count + 6'd1;
                end						  
					 6'd2:
					 begin
						  w16 <= (wt_16 ^ {wt_16[16:0],wt_16[31:17]} ^ {wt_16[8:0],wt_16[31:9]}) ^ {w3[24:0],w3[31:25]} ^ w10;
						  w17 <= (wt_17 ^ {wt_17[16:0],wt_17[31:17]} ^ {wt_17[8:0],wt_17[31:9]}) ^ {w4[24:0],w4[31:25]} ^ w11;
						  w18 <= (wt_18 ^ {wt_18[16:0],wt_18[31:17]} ^ {wt_18[8:0],wt_18[31:9]}) ^ {w5[24:0],w5[31:25]} ^ w12;
				        
						  count <= count + 6'd1;
					 end
					 6'd3:
					 begin
					     wt_19 <= w3 ^ w10 ^ {w16[16:0],w16[31:17]};
						  wt_20 <= w4 ^ w11 ^ {w17[16:0],w17[31:17]};
						  wt_21 <= w5 ^ w12 ^ {w18[16:0],w18[31:17]};
						  
						  w_12 <= w12 ^ w16;
						  w_13 <= w13 ^ w17;
						  w_14 <= w14 ^ w18;
						  
						  count <= count + 6'd1;
					 end
					 6'd4:
					 begin
					     w19 <= (wt_19 ^ {wt_19[16:0],wt_19[31:17]} ^ {wt_19[8:0],wt_19[31:9]}) ^ {w6[24:0],w6[31:25]} ^ w13;
						  w20 <= (wt_20 ^ {wt_20[16:0],wt_20[31:17]} ^ {wt_20[8:0],wt_20[31:9]}) ^ {w7[24:0],w7[31:25]} ^ w14;
						  w21 <= (wt_21 ^ {wt_21[16:0],wt_21[31:17]} ^ {wt_21[8:0],wt_21[31:9]}) ^ {w8[24:0],w8[31:25]} ^ w15;
					     
						  count <= count + 6'd1;
					 end
					 6'd5:
					 begin
					     wt_22 <= w6 ^ w13 ^ {w19[16:0],w19[31:17]};
						  wt_23 <= w7 ^ w14 ^ {w20[16:0],w20[31:17]};
						  wt_24 <= w8 ^ w15 ^ {w21[16:0],w21[31:17]};
						  
						  w_15 <= w15 ^ w19;
						  w_16 <= w16 ^ w20;
						  w_17 <= w17 ^ w21;
						  
						  count <= count + 6'd1;
					 end
					 6'd6:
					 begin
					     w22 <= (wt_22 ^ {wt_22[16:0],wt_22[31:17]} ^ {wt_22[8:0],wt_22[31:9]}) ^ {w9[24:0],w9[31:25]} ^ w16;
						  w23 <= (wt_23 ^ {wt_23[16:0],wt_23[31:17]} ^ {wt_23[8:0],wt_23[31:9]}) ^ {w10[24:0],w10[31:25]} ^ w17;
						  w24 <= (wt_24 ^ {wt_24[16:0],wt_24[31:17]} ^ {wt_24[8:0],wt_24[31:9]}) ^ {w11[24:0],w11[31:25]} ^ w18;	  
					 
					     count <= count + 6'd1;
					 end
					 6'd7:
					 begin
					     wt_25 <= w9 ^ w16 ^ {w22[16:0],w22[31:17]};
						  wt_26 <= w10 ^ w17 ^ {w23[16:0],w23[31:17]};
						  wt_27 <= w11 ^ w18 ^ {w24[16:0],w24[31:17]};
						  
						  w_18 <= w18 ^ w22;
						  w_19 <= w19 ^ w23;
						  w_20 <= w20 ^ w24;
						  
						  count <= count + 6'd1;
					 end
					 6'd8:
					 begin
					     w25 <= (wt_25 ^ {wt_25[16:0],wt_25[31:17]} ^ {wt_25[8:0],wt_25[31:9]}) ^ {w12[24:0],w12[31:25]} ^ w19;
						  w26 <= (wt_26 ^ {wt_26[16:0],wt_26[31:17]} ^ {wt_26[8:0],wt_26[31:9]}) ^ {w13[24:0],w13[31:25]} ^ w20;
						  w27 <= (wt_27 ^ {wt_27[16:0],wt_27[31:17]} ^ {wt_27[8:0],wt_27[31:9]}) ^ {w14[24:0],w14[31:25]} ^ w21;	  
					 
					     count <= count + 6'd1;
					 end
					 6'd9:
					 begin
					     wt_28 <= w12 ^ w19 ^ {w25[16:0],w25[31:17]};
						  wt_29 <= w13 ^ w20 ^ {w26[16:0],w26[31:17]};
						  wt_30 <= w14 ^ w21 ^ {w27[16:0],w27[31:17]};
						  
						  w_21 <= w21 ^ w25;
						  w_22 <= w22 ^ w26;
						  w_23 <= w23 ^ w27;
						  
						  count <= count + 6'd1;
					 end
					 6'd10:
					 begin
					     w28 <= (wt_28 ^ {wt_28[16:0],wt_28[31:17]} ^ {wt_28[8:0],wt_28[31:9]}) ^ {w15[24:0],w15[31:25]} ^ w22;
						  w29 <= (wt_29 ^ {wt_29[16:0],wt_29[31:17]} ^ {wt_29[8:0],wt_29[31:9]}) ^ {w16[24:0],w16[31:25]} ^ w23;
						  w30 <= (wt_30 ^ {wt_30[16:0],wt_30[31:17]} ^ {wt_30[8:0],wt_30[31:9]}) ^ {w17[24:0],w17[31:25]} ^ w24;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd11:
					 begin
					     wt_31 <= w15 ^ w22 ^ {w28[16:0],w28[31:17]};
						  wt_32 <= w16 ^ w23 ^ {w29[16:0],w29[31:17]};
						  wt_33 <= w17 ^ w24 ^ {w30[16:0],w30[31:17]};
						  
						  w_24 <= w24 ^ w28;
						  w_25 <= w25 ^ w29;
						  w_26 <= w26 ^ w30;
						  
						  count <= count + 6'd1;
					 end
					 6'd12:
					 begin
					     w31 <= (wt_31 ^ {wt_31[16:0],wt_31[31:17]} ^ {wt_31[8:0],wt_31[31:9]}) ^ {w18[24:0],w18[31:25]} ^ w25;
						  w32 <= (wt_32 ^ {wt_32[16:0],wt_32[31:17]} ^ {wt_32[8:0],wt_32[31:9]}) ^ {w19[24:0],w19[31:25]} ^ w26;
						  w33 <= (wt_33 ^ {wt_33[16:0],wt_33[31:17]} ^ {wt_33[8:0],wt_33[31:9]}) ^ {w20[24:0],w20[31:25]} ^ w27;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd13:
					 begin
					     wt_34 <= w18 ^ w25 ^ {w31[16:0],w31[31:17]};
						  wt_35 <= w19 ^ w26 ^ {w32[16:0],w32[31:17]};
						  wt_36 <= w20 ^ w27 ^ {w33[16:0],w33[31:17]};
						  
						  w_27 <= w27 ^ w31;
						  w_28 <= w28 ^ w32;
						  w_29 <= w29 ^ w33;
						  
						  count <= count + 6'd1;
					 end
					 6'd14:
					 begin
					     w34 <= (wt_34 ^ {wt_34[16:0],wt_34[31:17]} ^ {wt_34[8:0],wt_34[31:9]}) ^ {w21[24:0],w21[31:25]} ^ w28;
						  w35 <= (wt_35 ^ {wt_35[16:0],wt_35[31:17]} ^ {wt_35[8:0],wt_35[31:9]}) ^ {w22[24:0],w22[31:25]} ^ w29;
						  w36 <= (wt_36 ^ {wt_36[16:0],wt_36[31:17]} ^ {wt_36[8:0],wt_36[31:9]}) ^ {w23[24:0],w23[31:25]} ^ w30;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd15:
					 begin
					     wt_37 <= w21 ^ w28 ^ {w34[16:0],w34[31:17]};
						  wt_38 <= w22 ^ w29 ^ {w35[16:0],w35[31:17]};
						  wt_39 <= w23 ^ w30 ^ {w36[16:0],w36[31:17]};
						  
						  w_30 <= w30 ^ w34;
						  w_31 <= w31 ^ w35;
						  w_32 <= w32 ^ w36;
						  
						  count <= count + 6'd1;
					 end
					 6'd16:
					 begin
					     w37 <= (wt_37 ^ {wt_37[16:0],wt_37[31:17]} ^ {wt_37[8:0],wt_37[31:9]}) ^ {w24[24:0],w24[31:25]} ^ w31;
						  w38 <= (wt_38 ^ {wt_38[16:0],wt_38[31:17]} ^ {wt_38[8:0],wt_38[31:9]}) ^ {w25[24:0],w25[31:25]} ^ w32;
						  w39 <= (wt_39 ^ {wt_39[16:0],wt_39[31:17]} ^ {wt_39[8:0],wt_39[31:9]}) ^ {w26[24:0],w26[31:25]} ^ w33;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd17:
					 begin
					     wt_40 <= w24 ^ w31 ^ {w37[16:0],w37[31:17]};
						  wt_41 <= w25 ^ w32 ^ {w38[16:0],w38[31:17]};
						  wt_42 <= w26 ^ w33 ^ {w39[16:0],w39[31:17]};
						  
						  w_33 <= w33 ^ w37;
						  w_34 <= w34 ^ w38;
						  w_35 <= w35 ^ w39;
						  
						  count <= count + 6'd1;
					 end
					 6'd18:
					 begin
					     w40 <= (wt_40 ^ {wt_40[16:0],wt_40[31:17]} ^ {wt_40[8:0],wt_40[31:9]}) ^ {w27[24:0],w27[31:25]} ^ w34;
						  w41 <= (wt_41 ^ {wt_41[16:0],wt_41[31:17]} ^ {wt_41[8:0],wt_41[31:9]}) ^ {w28[24:0],w28[31:25]} ^ w35;
						  w42 <= (wt_42 ^ {wt_42[16:0],wt_42[31:17]} ^ {wt_42[8:0],wt_42[31:9]}) ^ {w29[24:0],w29[31:25]} ^ w36;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd19:
					 begin
					     wt_43 <= w27 ^ w34 ^ {w40[16:0],w40[31:17]};
						  wt_44 <= w28 ^ w35 ^ {w41[16:0],w41[31:17]};
						  wt_45 <= w29 ^ w36 ^ {w42[16:0],w42[31:17]};
						  
						  w_36 <= w36 ^ w40;
						  w_37 <= w37 ^ w41;
						  w_38 <= w38 ^ w42;
						  
						  count <= count + 6'd1;
					 end
					 6'd20:
					 begin
					     w43 <= (wt_43 ^ {wt_43[16:0],wt_43[31:17]} ^ {wt_43[8:0],wt_43[31:9]}) ^ {w30[24:0],w30[31:25]} ^ w37;
						  w44 <= (wt_44 ^ {wt_44[16:0],wt_44[31:17]} ^ {wt_44[8:0],wt_44[31:9]}) ^ {w31[24:0],w31[31:25]} ^ w38;
						  w45 <= (wt_45 ^ {wt_45[16:0],wt_45[31:17]} ^ {wt_45[8:0],wt_45[31:9]}) ^ {w32[24:0],w32[31:25]} ^ w39;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd21:
					 begin
					     wt_46 <= w30 ^ w37 ^ {w43[16:0],w43[31:17]};
						  wt_47 <= w31 ^ w38 ^ {w44[16:0],w44[31:17]};
						  wt_48 <= w32 ^ w39 ^ {w45[16:0],w45[31:17]};
						  
						  w_39 <= w39 ^ w43;
						  w_40 <= w40 ^ w44;
						  w_41 <= w41 ^ w45;
						  
						  count <= count + 6'd1;
					 end
					 6'd22:
					 begin
					     w46 <= (wt_46 ^ {wt_46[16:0],wt_46[31:17]} ^ {wt_46[8:0],wt_46[31:9]}) ^ {w33[24:0],w33[31:25]} ^ w40;
						  w47 <= (wt_47 ^ {wt_47[16:0],wt_47[31:17]} ^ {wt_47[8:0],wt_47[31:9]}) ^ {w34[24:0],w34[31:25]} ^ w41;
						  w48 <= (wt_48 ^ {wt_48[16:0],wt_48[31:17]} ^ {wt_48[8:0],wt_48[31:9]}) ^ {w35[24:0],w35[31:25]} ^ w42;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd23:
					 begin
					     wt_49 <= w33 ^ w40 ^ {w46[16:0],w46[31:17]};
						  wt_50 <= w34 ^ w41 ^ {w47[16:0],w47[31:17]};
						  wt_51 <= w35 ^ w42 ^ {w48[16:0],w48[31:17]};
						  
						  w_42 <= w42 ^ w46;
						  w_43 <= w43 ^ w47;
						  w_44 <= w44 ^ w48;
						  
						  count <= count + 6'd1;
					 end
					 6'd24:
					 begin
					     w49 <= (wt_49 ^ {wt_49[16:0],wt_49[31:17]} ^ {wt_49[8:0],wt_49[31:9]}) ^ {w36[24:0],w36[31:25]} ^ w43;
						  w50 <= (wt_50 ^ {wt_50[16:0],wt_50[31:17]} ^ {wt_50[8:0],wt_50[31:9]}) ^ {w37[24:0],w37[31:25]} ^ w44;
						  w51 <= (wt_51 ^ {wt_51[16:0],wt_51[31:17]} ^ {wt_51[8:0],wt_51[31:9]}) ^ {w38[24:0],w38[31:25]} ^ w45;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd25:
					 begin
					     wt_52 <= w36 ^ w43 ^ {w49[16:0],w49[31:17]};
						  wt_53 <= w37 ^ w44 ^ {w50[16:0],w50[31:17]};
						  wt_54 <= w38 ^ w45 ^ {w51[16:0],w51[31:17]};
						  
						  w_45 <= w45 ^ w49;
						  w_46 <= w46 ^ w50;
						  w_47 <= w47 ^ w51;
						  
						  count <= count + 6'd1;
					 end
					 6'd26:
					 begin
					     w52 <= (wt_52 ^ {wt_52[16:0],wt_52[31:17]} ^ {wt_52[8:0],wt_52[31:9]}) ^ {w39[24:0],w39[31:25]} ^ w46;
						  w53 <= (wt_53 ^ {wt_53[16:0],wt_53[31:17]} ^ {wt_53[8:0],wt_53[31:9]}) ^ {w40[24:0],w40[31:25]} ^ w47;
						  w54 <= (wt_54 ^ {wt_54[16:0],wt_54[31:17]} ^ {wt_54[8:0],wt_54[31:9]}) ^ {w41[24:0],w41[31:25]} ^ w48;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd27:
					 begin
					     wt_55 <= w39 ^ w46 ^ {w52[16:0],w52[31:17]};
						  wt_56 <= w40 ^ w47 ^ {w53[16:0],w53[31:17]};
						  wt_57 <= w41 ^ w48 ^ {w54[16:0],w54[31:17]};
						  
						  w_48 <= w48 ^ w52;
						  w_49 <= w49 ^ w53;
						  w_50 <= w50 ^ w54;
						  
						  count <= count + 6'd1;
					 end
					 6'd28:
					 begin
					     w55 <= (wt_55 ^ {wt_55[16:0],wt_55[31:17]} ^ {wt_55[8:0],wt_55[31:9]}) ^ {w42[24:0],w42[31:25]} ^ w49;
						  w56 <= (wt_56 ^ {wt_56[16:0],wt_56[31:17]} ^ {wt_56[8:0],wt_56[31:9]}) ^ {w43[24:0],w43[31:25]} ^ w50;
						  w57 <= (wt_57 ^ {wt_57[16:0],wt_57[31:17]} ^ {wt_57[8:0],wt_57[31:9]}) ^ {w44[24:0],w44[31:25]} ^ w51;	  
					 
					     count <= count + 6'd1;
					 end
			       6'd29:
					 begin
					     wt_58 <= w42 ^ w49 ^ {w55[16:0],w55[31:17]};
						  wt_59 <= w43 ^ w50 ^ {w56[16:0],w56[31:17]};
						  wt_60 <= w44 ^ w51 ^ {w57[16:0],w57[31:17]};
						  
						  w_51 <= w51 ^ w55;
						  w_52 <= w52 ^ w56;
						  w_53 <= w53 ^ w57;
						  
						  count <= count + 6'd1;
					 end
					 6'd30:
					 begin
					     w58 <= (wt_58 ^ {wt_58[16:0],wt_58[31:17]} ^ {wt_58[8:0],wt_58[31:9]}) ^ {w45[24:0],w45[31:25]} ^ w52;
						  w59 <= (wt_59 ^ {wt_59[16:0],wt_59[31:17]} ^ {wt_59[8:0],wt_59[31:9]}) ^ {w46[24:0],w46[31:25]} ^ w53;
						  w60 <= (wt_60 ^ {wt_60[16:0],wt_60[31:17]} ^ {wt_60[8:0],wt_60[31:9]}) ^ {w47[24:0],w47[31:25]} ^ w54;	  
					 
					     count <= count + 6'd1;
					 end		
					 6'd31:
					 begin
					     wt_61 <= w45 ^ w52 ^ {w58[16:0],w58[31:17]};
						  wt_62 <= w46 ^ w53 ^ {w59[16:0],w59[31:17]};
						  wt_63 <= w47 ^ w54 ^ {w60[16:0],w60[31:17]};
						  
						  w_54 <= w54 ^ w58;
						  w_55 <= w55 ^ w59;
						  w_56 <= w56 ^ w60;
						  
						  count <= count + 6'd1;
					 end
					 6'd32:
					 begin
					     w61 <= (wt_61 ^ {wt_61[16:0],wt_61[31:17]} ^ {wt_61[8:0],wt_61[31:9]}) ^ {w48[24:0],w48[31:25]} ^ w55;
						  w62 <= (wt_62 ^ {wt_62[16:0],wt_62[31:17]} ^ {wt_62[8:0],wt_62[31:9]}) ^ {w49[24:0],w49[31:25]} ^ w56;
						  w63 <= (wt_63 ^ {wt_63[16:0],wt_63[31:17]} ^ {wt_63[8:0],wt_63[31:9]}) ^ {w50[24:0],w50[31:25]} ^ w57;	  
					 
					     count <= count + 6'd1;
					 end
					 6'd33:
					 begin
					     wt_64 <= w48 ^ w55 ^ {w61[16:0],w61[31:17]};
						  wt_65 <= w49 ^ w56 ^ {w62[16:0],w62[31:17]};
						  wt_66 <= w50 ^ w57 ^ {w63[16:0],w63[31:17]};
						  
						  w_57 <= w57 ^ w61;
						  w_58 <= w58 ^ w62;
						  w_59 <= w59 ^ w63;
						  
						  count <= count + 6'd1;
					 end
					 6'd34:
					 begin
					     w64 <= (wt_64 ^ {wt_64[16:0],wt_64[31:17]} ^ {wt_64[8:0],wt_64[31:9]}) ^ {w51[24:0],w51[31:25]} ^ w58;
						  w65 <= (wt_65 ^ {wt_65[16:0],wt_65[31:17]} ^ {wt_65[8:0],wt_65[31:9]}) ^ {w52[24:0],w52[31:25]} ^ w59;
						  w66 <= (wt_66 ^ {wt_66[16:0],wt_66[31:17]} ^ {wt_66[8:0],wt_66[31:9]}) ^ {w53[24:0],w53[31:25]} ^ w60;	  
					 
					     count <= count + 6'd1;
					 end
					 6'd35:
					 begin
					     wt_67 <= w51 ^ w58 ^ {w64[16:0],w64[31:17]};
						  
						  w_60 <= w60 ^ w64;
						  w_61 <= w61 ^ w65;
						  w_62 <= w62 ^ w66;
						  						  
						  count <= count + 6'd1;
					 end
					 6'd36:
					 begin
					     w67 <= (wt_67 ^ {wt_67[16:0],wt_67[31:17]} ^ {wt_67[8:0],wt_67[31:9]}) ^ {w54[24:0],w54[31:25]} ^ w61;
					     
						  count <= count + 6'd1;
					 end
                6'd37:
					 begin
					     w_63 <= w63 ^ w67;
						  
					     count <= 6'd0;//清零
					 end
					 
					 default:
					 begin
					     count <= 6'd0;
					 end
				endcase
		  end
	 end
	 

	 
	 
/*
    always@(posedge clk or negedge rst)
    begin
        if(!rst)
		  begin
		      Tj <= 32'h79CC4519;
				FF <= A ^ B ^ C;
				GG <= E ^ F ^ G;
		  end
		  else if(!enable)
		  begin
		      Tj <= Tj;
				FF <= FF;
				GG <= GG;
		  end
		  else if(j >= 6'd15 && j<= 6'd62)
		  begin
      		Tj <= 32'h7A879D8A;
				FF <= ((A & B) | (B & C) | (A & C) );
				GG <= ((E & F) | (~E & G));				
		  end
		  else
		  begin
		      
            Tj <= 32'h79CC4519;
				FF <= A ^ B ^ C;
				GG <= E ^ F ^ G;				
		  end
    end
*/	 
	
	 
	 always@(posedge clk or negedge rst)
	 begin
	     if(!rst)
		  begin
		      V_o <= 256'd0;       //复位时回归默认值
				j <= 6'd0;
				{A,B,C,D,E,F,G,H} <= 256'd0;
				
				Tj <= 32'h79CC4519;
				FF <= A ^ B ^ C;
				GG <= E ^ F ^ G;
		  end
		  else if(!enable)
		  begin       
		      V_o <= V_o;          //使能无效时暂停工作
				j <= j;
				{A,B,C,D,E,F,G,H} <= {A,B,C,D,E,F,G,H};
				
				Tj <= Tj;
				FF <= FF;
				GG <= GG;
		  end
		  else 
		  begin
		      case(j)
				    6'd0:
					 begin
					     {A,B,C,D,E,F,G,H} = V_i;//寄存器赋初值
							
					     if(count == 6'd2)//判断w0与w_0是否已计算完成
						  begin
						      Tj = 32'h79CC4519;//完成则开始第一次逻辑运算
				            FF = A ^ B ^ C;
				            GG = E ^ F ^ G;
								
						      SS1t = {A[19:0],A[31:20]} + E + Tj;
							   SS1 = {SS1t[24:0],SS1t[31:25]};
							   SS2 = SS1 ^ {A[19:0],A[31:20]};
							   TT1 = FF + D + SS2 + w_0;
							   TT2 = GG + H + SS1 + w0;
							
							   D = C;
							   C = {B[22:0],B[31:23]};
							   B = A;
							   A = TT1;
							   H = G;
							   G = {F[12:0],F[31:13]};
							   F = E;
							   E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};
							
							   j = j + 6'd1;
						  end
						  else
						  begin
						      j = j;//未完成则保持j不变，下一个clk重复判断
					     end
					 end
				    6'd1:
					 begin
					     Tj = 32'h79CC4519;//第二次逻辑运算
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
								
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[30:0],Tj[31]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_1;
						  TT2 = GG + H + SS1 + w1;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};
						  
						  j = j + 6'd1;
					 end
		          6'd2:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[29:0],Tj[31:30]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_2;
						  TT2 = GG + H + SS1 + w2;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};
						  
						  j = j + 6'd1;
					 end
					 6'd3:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[28:0],Tj[31:29]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_3;
						  TT2 = GG + H + SS1 + w3;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd4:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[27:0],Tj[31:28]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_4;
						  TT2 = GG + H + SS1 + w4;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd5:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[26:0],Tj[31:27]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_5;
						  TT2 = GG + H + SS1 + w5;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd6:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[25:0],Tj[31:26]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_6;
						  TT2 = GG + H + SS1 + w6;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd7:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[24:0],Tj[31:25]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_7;
						  TT2 = GG + H + SS1 + w7;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd8:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[23:0],Tj[31:24]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_8;
						  TT2 = GG + H + SS1 + w8;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd9:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[22:0],Tj[31:23]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_9;
						  TT2 = GG + H + SS1 + w9;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd10:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[21:0],Tj[31:22]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_10;
						  TT2 = GG + H + SS1 + w10;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};
						  
					     j = j + 6'd1;
					 end
					 6'd11:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[20:0],Tj[31:21]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_11;
						  TT2 = GG + H + SS1 + w11;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};
						  
					     j = j + 6'd1;
					 end
					 6'd12:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[19:0],Tj[31:20]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_12;
						  TT2 = GG + H + SS1 + w12;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd13:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[18:0],Tj[31:19]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_13;
						  TT2 = GG + H + SS1 + w13;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};	     
						  
					     j = j + 6'd1;
					 end
					 6'd14:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[17:0],Tj[31:18]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_14;
						  TT2 = GG + H + SS1 + w14;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd15:
					 begin
					     Tj = 32'h79CC4519;
				        FF = A ^ B ^ C;
				        GG = E ^ F ^ G;
							
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[16:0],Tj[31:17]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_15;
						  TT2 = GG + H + SS1 + w15;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd16:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[15:0],Tj[31:16]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_16;
						  TT2 = GG + H + SS1 + w16;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd17:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[14:0],Tj[31:15]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_17;
						  TT2 = GG + H + SS1 + w17;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};		     
						  
					     j = j + 6'd1;
					 end
					 6'd18:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[13:0],Tj[31:14]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_18;
						  TT2 = GG + H + SS1 + w18;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};     
						  
					     j = j + 6'd1;
					 end
					 6'd19:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[12:0],Tj[31:13]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_19;
						  TT2 = GG + H + SS1 + w19;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};	     
						  
					     j = j + 6'd1;
					 end
					 6'd20:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[11:0],Tj[31:12]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_20;
						  TT2 = GG + H + SS1 + w20;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};     
						  
					     j = j + 6'd1;
					 end
					 6'd21:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[10:0],Tj[31:11]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_21;
						  TT2 = GG + H + SS1 + w21;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};		     
						  
					     j = j + 6'd1;
					 end
					 6'd22:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[9:0],Tj[31:10]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_22;
						  TT2 = GG + H + SS1 + w22;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};     
						  
					     j = j + 6'd1;
					 end
					 6'd23:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[8:0],Tj[31:9]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_23;
						  TT2 = GG + H + SS1 + w23;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};	     
						  
					     j = j + 6'd1;
					 end
					 6'd24:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[7:0],Tj[31:8]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_24;
						  TT2 = GG + H + SS1 + w24;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd25:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[6:0],Tj[31:7]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_25;
						  TT2 = GG + H + SS1 + w25;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};		     
						  
					     j = j + 6'd1;
					 end
					 6'd26:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[5:0],Tj[31:6]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_26;
						  TT2 = GG + H + SS1 + w26;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd27:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[4:0],Tj[31:5]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_27;
						  TT2 = GG + H + SS1 + w27;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd28:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[3:0],Tj[31:4]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_28;
						  TT2 = GG + H + SS1 + w28;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd29:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[2:0],Tj[31:3]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_29;
						  TT2 = GG + H + SS1 + w29;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd30:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[1:0],Tj[31:2]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_30;
						  TT2 = GG + H + SS1 + w30;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd31:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[0],Tj[31:1]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_31;
						  TT2 = GG + H + SS1 + w31;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd32:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + Tj;
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_32;
						  TT2 = GG + H + SS1 + w32;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd33:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[30:0],Tj[31]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_33;
						  TT2 = GG + H + SS1 + w33;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd34:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[29:0],Tj[31:30]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_34;
						  TT2 = GG + H + SS1 + w34;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd35:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[28:0],Tj[31:29]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_35;
						  TT2 = GG + H + SS1 + w35;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd36:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[27:0],Tj[31:28]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_36;
						  TT2 = GG + H + SS1 + w36;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd37:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[26:0],Tj[31:27]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_37;
						  TT2 = GG + H + SS1 + w37;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd38:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[25:0],Tj[31:26]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_38;
						  TT2 = GG + H + SS1 + w38;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd39:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[24:0],Tj[31:25]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_39;
						  TT2 = GG + H + SS1 + w39;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd40:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[23:0],Tj[31:24]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_40;
						  TT2 = GG + H + SS1 + w40;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd41:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[22:0],Tj[31:23]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_41;
						  TT2 = GG + H + SS1 + w41;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd42:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[21:0],Tj[31:22]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_42;
						  TT2 = GG + H + SS1 + w42;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd43:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[20:0],Tj[31:21]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_43;
						  TT2 = GG + H + SS1 + w43;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd44:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[19:0],Tj[31:20]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_44;
						  TT2 = GG + H + SS1 + w44;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd45:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[18:0],Tj[31:19]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_45;
						  TT2 = GG + H + SS1 + w45;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd46:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[17:0],Tj[31:18]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_46;
						  TT2 = GG + H + SS1 + w46;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd47:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[16:0],Tj[31:17]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_47;
						  TT2 = GG + H + SS1 + w47;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd48:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[15:0],Tj[31:16]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_48;
						  TT2 = GG + H + SS1 + w48;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd49:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[14:0],Tj[31:15]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_49;
						  TT2 = GG + H + SS1 + w49;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd50:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[13:0],Tj[31:14]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_50;
						  TT2 = GG + H + SS1 + w50;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd51:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[12:0],Tj[31:13]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_51;
						  TT2 = GG + H + SS1 + w51;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd52:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[11:0],Tj[31:12]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_52;
						  TT2 = GG + H + SS1 + w52;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd53:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[10:0],Tj[31:11]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_53;
						  TT2 = GG + H + SS1 + w53;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd54:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[9:0],Tj[31:10]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_54;
						  TT2 = GG + H + SS1 + w54;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};			     
						  
					     j = j + 6'd1;
					 end
					 6'd55:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[8:0],Tj[31:9]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_55;
						  TT2 = GG + H + SS1 + w55;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd56:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[7:0],Tj[31:8]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_56;
						  TT2 = GG + H + SS1 + w56;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd57:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[6:0],Tj[31:7]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_57;
						  TT2 = GG + H + SS1 + w57;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd58:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[5:0],Tj[31:6]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_58;
						  TT2 = GG + H + SS1 + w58;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd59:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[4:0],Tj[31:5]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_59;
						  TT2 = GG + H + SS1 + w59;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd60:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[3:0],Tj[31:4]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_60;
						  TT2 = GG + H + SS1 + w60;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};					     
						  
					     j = j + 6'd1;
					 end
					 6'd61:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[2:0],Tj[31:3]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_61;
						  TT2 = GG + H + SS1 + w61;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd62:
					 begin
		              Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[1:0],Tj[31:2]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_62;
						  TT2 = GG + H + SS1 + w62;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
					     j = j + 6'd1;
					 end
					 6'd63:
					 begin
					     Tj = 32'h7A879D8A;
				        FF = ((A & B) | (B & C) | (A & C) );
				        GG = ((E & F) | (~E & G));	
						  
					     SS1t = {A[19:0],A[31:20]} + E + {Tj[0],Tj[31:1]};
						  SS1 = {SS1t[24:0],SS1t[31:25]};
						  SS2 = SS1 ^ {A[19:0],A[31:20]};
						  TT1 = FF + D + SS2 + w_63;
						  TT2 = GG + H + SS1 + w63;
							
						  D = C;
						  C = {B[22:0],B[31:23]};
						  B = A;
						  A = TT1;
						  H = G;
						  G = {F[12:0],F[31:13]};
						  F = E;
						  E = TT2 ^ {TT2[22:0],TT2[31:23]} ^ {TT2[14:0],TT2[31:15]};				     
						  
						  V_o = {A,B,C,D,E,F,G,H} ^ V_i;//输出
						  
					     j = 6'd0;//64次逻辑运算完成后回归初态
					 end
					 default:
					 begin
					     j = 6'd0;
					 end
				endcase
		  end
	 end
	 
endmodule
